﻿* Transient Analysis, 4.2E3 bandPass, 4th order Chebyshev undefined dB, 2 stages using AD8542

* Input signal for AC and Transient (step) analysis 
VIN IN 0 AC 1 DC 2.5 PULSE(2.5 4.89 0ns 1ns 1ns 1s 2s) 
* VNOISE IN 0 AC 0 DC 2.5 

XA IN OUTA VCCG VEEG VREF sallenKeylowPassStageA
XB OUTA OUT VCCG VEEG VREF sallenKeyhighPassStageB

VP VCCG 0 5
VM VEEG 0 0
VR VREF 0 2.5

*Simulation directive lines for Transient Analysis 
.TRAN 1ns 1.5E-3 
*.AC DEC 100 11.3 80E3 
*.NOISE V(OUT) VNOISE DEC 100 11.3 80E3 
.PROBE 

.SUBCKT sallenKeylowPassStageA IN OUT VCC VEE REF 
X1 INP OUT VCC VEE OUT  AD8542 
R1 IN 1  8.45E3 
R2 1 INP 118E3 
C1 1 OUT 3.9E-9 
C2 INP REF 390E-12 
.ENDS sallenKeylowPassStageA 

.SUBCKT sallenKeyhighPassStageB IN OUT VCC VEE REF 
X1 INP OUT VCC VEE OUT  AD8542 
C1 IN 1 68E-9 
C2 1 INP 68E-9 
R1 1 OUT  6.34E3 
R2 INP REF 15.8E3 
.ENDS sallenKeyhighPassStageB 

* AD8542 SPICE Macro-model Typical Values
* Description: Amplifier
* Generic Desc: 2.7/5V, CMOS, OP, Low Pwr, RRIO, 2X
* Developed by: TAM / ADSC
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (06/1998)
* Copyright 1998, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node Assignments
*		noninverting input
*		|	inverting input
*		|	|	 positive supply
*		|	|	 |	 negative supply
*		|	|	 |	 |	 output
*		|	|	 |	 |	 |
*		|	|	 |	 |	 |
.SUBCKT AD8542	1	2	99	50	45
*
* INPUT STAGE
*
M1   4  1 8 8 PIX L=0.6E-6 W=16E-6
M2   6  7 8 8 PIX L=0.6E-6 W=16E-6
M3  11  1 10 10 NIX L=0.6E-6 W=16E-6
M4  12  7 10 10 NIX L=0.6E-6 W=16E-6
RC1  4 50 20E3
RC2  6 50 20E3
RC3 99 11 20E3
RC4 99 12 20E3
C1   4  6 1.5E-12
C2  11 12 1.5E-12
I1  99  8 1E-5
I2  10 50 1E-5
V1  99  9 0.2
V2  13 50 0.2
D1   8  9 DX
D2  13 10 DX
EOS  7  2 POLY(3) (22,98) (73,98) (81,0) 1E-3 1 1 1
IOS  1  2 2.5E-12
*
* CMRR 64dB, ZERO AT 20kHz
*
ECM1 21 98 POLY(2) (1,98) (2,98) 0 .5 .5
RCM1 21 22 79.6E3
CCM1 21 22 100E-12
RCM2 22 98 50
*
* PSRR=90dB, ZERO AT 200Hz
*
RPS1 70  0 1E6
RPS2 71  0 1E6
CPS1 99 70 1E-5
CPS2 50 71 1E-5
EPSY 98 72 POLY(2) (70,0) (0,71) 0 1 1
RPS3 72 73 1.59E6
CPS3 72 73 500E-12
RPS4 73 98 25
*
* VOLTAGE NOISE REFERENCE OF 35nV/rt(Hz)
*
VN1 80 0 0
RN1 80 0 16.45E-3
HN  81 0 VN1 35
RN2 81 0 1
*
* INTERNAL VOLTAGE REFERENCE
*
VFIX 90 98 DC 1
S1   90 91 (50,99) VSY_SWITCH
VSN1 91 92 DC 0
RSY  92 98 1E3
EREF 98  0 POLY(2) (99,0) (50,0) 0 .5 .5
GSY  99 50 POLY(1) (99,50) 0 3.7E-6
*
* ADAPTIVE GAIN STAGE
* AT Vsy>+4.2, AVol=45  V/mv
* AT Vsy<+3.8, AVol=450 V/mv
*
G1  98 30 POLY(2) (4,6) (11,12) 0 2.5E-5 2.5E-5
VR1 30 31 DC 0
H1  31 98 POLY(2) VR1 VSN1 0 5.45E6 0 0 49.05E9
CF  45 30 10E-12
D3  30 99 DX
D4  50 30 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=0.6E-6 W=375E-6
M6  45 47 50 50 NOX L=0.6E-6 W=500E-6
EG1 99 46 POLY(1) (98,30) 1.05 1
EG2 47 50 POLY(1) (30,98) 1.04 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=20E-6,VTO=-1,LAMBDA=0.067)
.MODEL NOX NMOS (LEVEL=2,KP=20E-6,VTO=1,LAMBDA=0.067)
.MODEL PIX PMOS (LEVEL=2,KP=20E-6,VTO=-0.7,LAMBDA=0.01,KF=1E-31)
.MODEL NIX NMOS (LEVEL=2,KP=20E-6,VTO=0.7,LAMBDA=0.01,KF=1E-31)
.MODEL DX D(IS=1E-14)
.MODEL VSY_SWITCH VSWITCH(ROFF=100E3,RON=1,VOFF=-4.2,VON=-3.5)
.ENDS AD8542




